`ifndef MIPS_H
`include "mips.h"
`endif

`ifndef EXECUTE_STAGE
`define EXECUTE_STAGE

`include "execute/alu.v"
`include "execute/execute_pipeline_reg.v"
`include "util.v"

// This module encapsulates the entire execute stage.
module execute_stage(clk, FlushE, RegWriteD, MemtoRegD, MemWriteD, ALUControlD,
	ALUSrcD, RegDstD, RD1D, RD2D, RsD, RtD, RdD, SignImmD,
	RegWriteE, MemtoRegE, MemWriteE, RegDstE, ALUControlE,
	RD1E, RD2E, RsE, RtE, RdE, SignImmE, shamtD, 
	ResultW, ALUOutM, ForwardAE, ForwardBE,
	WriteRegE, WriteDataE, ALUOutE);

	// The clock.
	input wire clk;

	// The flag from the Hazard Unit raised when this pipeline stage should be
	// flushed.
	input wire FlushE;

	/*** The following inputs are fed from the Decode pipeline stage ***/

	// The control signal denoting whether a register is written to.
	input wire RegWriteD;

	// The control signal denoting whether data is being written from
	// memory to a register.
	input wire MemtoRegD;

	// The control signal denoting whether main memory is being written to.
	input wire MemWriteD;

	// The four-bit ALU op denoting which operation the ALU should perform.
	input wire [3:0] ALUControlD;

	// The control signal denoting whether the ALU input is an immediate value.
	input wire ALUSrcD;

	// The control signal denoting whether the write reg is rd (R-type instr).
	input wire RegDstD;

	// The data read from the first source register (rs).
	input wire [31:0] RD1D;

	// The data read from the second source register (rt).
	input wire [31:0] RD2D;

	// The first source register.
	input wire [4:0] RsD;

	// The second source register.
	input wire [4:0] RtD;

	// The destination register.
	input wire [4:0] RdD;

	// The sign-extended immediate value.
	input wire [31:0] SignImmD;

	/*** The following inputs are fed from elsewhere ***/

	// The chosen value to write (may be ALU output or from data memory).
	input wire [31:0] ResultW;

	// The output of the ALU after it has passed through the Memory pipeline reg.
	input wire [31:0] ALUOutM;

	// The input to the mux (from Hazard Unit) that determines SrcAE.
	input wire [1:0] ForwardAE;

	// The input to the mux (from Hazard Unit) that determines SrcBE.
	input wire [1:0] ForwardBE;

	/*** The following outputs are generated by the Execute pipeline stage ***/

	// The control signal denoting whether a register is written to.
	output wire RegWriteE;

	// The control signal denoting whether data is being written from
	// memory to a register.
	output wire MemtoRegE;

	// The control signal denoting whether main memory is being written to.
	output wire MemWriteE;

	// The four-bit ALU op denoting which operation the ALU should perform.
	output wire [3:0] ALUControlE;

	// The control signal denoting whether the ALU input is an immediate value.
	wire ALUSrcE;

	// The control signal denoting whether the write reg is rd (R-type instr).
	output wire RegDstE;

	// The data read from the first source register (rs).
	output wire [31:0] RD1E;

	// The data read from the second source register (rt).
	output wire [31:0] RD2E;

	// The first source register.
	output wire [4:0] RsE;

	// The second source register.
	output wire [4:0] RtE;

	// The destination register.
	output wire [4:0] RdE;

	// The sign-extended immediate value.
	output wire [31:0] SignImmE;

    // The shift amount value
    input wire [4:0] shamtD;
	/*** The following outputs are generated internal to the execute stage ***/

	// The 5-bit register code that will be written to.
	output wire [4:0] WriteRegE;

	// The 32-bit data to write to memory.
	output wire [31:0] WriteDataE;

	// The 32-bit LHS of the ALU operation to perform.
	wire [31:0] SrcAE; // Note: Not a top-level output from the EX stage

	// The 32-bit RHS of the ALU operation to perform.
	wire [31:0] SrcBE; // Note: Not a top-level output from the EX stage

    // The execute stage's shift immediate value
    wire [4:0] shamtE;

	// The 32-bit output from the ALU.
	output wire [31:0] ALUOutE;

	// Instantiate all muxes, the ALU, and the EX pipeline register

	execute_pipeline_reg EX_pipeline_reg(clk, FlushE, RegWriteD, MemtoRegD, MemWriteD,
		ALUControlD, ALUSrcD, RegDstD, RD1D, RD2D, RsD, RtD, RdD, SignImmD, shamtD
		RegWriteE, MemtoRegE, MemWriteE, ALUControlE, ALUSrcE, RegDstE,
		RD1E, RD2E, RsE, RtE, RdE, SignImmE, shamtE);

	mux5_2 write_reg_mux(RdE, RtE, RegDstE, WriteRegE);
	mux32_3 write_data_mux(RD2E, ResultW, ALUOutM, ForwardBE, WriteDataE);
	mux32_3 srcA_mux(RD1E, ResultW, ALUOutM, ForwardAE, SrcAE);
	mux32_2 srcB_mux(SignImmE, WriteDataE, ALUSrcE, SrcBE);

	alu myALU(SrcAE, SrcBE, ALUControlE, shamtE, ALUOutE);

endmodule
`endif

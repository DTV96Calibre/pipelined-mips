`ifndef MIPS_H
`include "mips.h"
`endif

`ifndef EXECUTE_PIPELINE_REG
`define EXECUTE_PIPELINE_REG

`include "register/pipeline_reg.v"

// This module encapsulates the entire execute pipeline register.
module execute_pipeline_reg(clk, FlushE, RegWriteD, MemtoRegD, MemWriteD, ALUControlD,
	ALUSrcD, RegDstD, RD1D, RD2D, RsD, RtD, RdD, SignImmD,
	RegWriteE, MemtoRegE, MemWriteE, ALUControlE, ALUSrcE, RegDstE,
	RD1E, RD2E, RsE, RtE, RdE, SignImmE);

	// The clock.
	input wire clk;

	// The flag from the Hazard Unit raised when this pipeline stage should be
	// flushed.
	input wire FlushE;

	/*** The following inputs are fed from the Decode pipeline stage ***/

	// The control signal denoting whether a register is written to.
	input wire RegWriteD;

	// The control signal denoting whether data is being written from
	// memory to a register.
	input wire MemtoRegD;

	// The control signal denoting whether main memory is being written to.
	input wire MemWriteD;

	// The four-bit ALU op denoting which operation the ALU should perform.
	input wire [3:0] ALUControlD;

	// The control signal denoting whether the ALU input is an immediate value.
	input wire ALUSrcD;

	// The control signal denoting whether the write reg is rd (R-type instr).
	input wire RegDstD;

	// The data read from the first source register (rs).
	input wire [31:0] RD1D;

	// The data read from the second source register (rt).
	input wire [31:0] RD2D;

	// The first source register.
	input wire [4:0] RsD;

	// The second source register.
	input wire [4:0] RtD;

	// The destination register.
	input wire [4:0] RdD;

	// The sign-extended immediate value.
	input wire [31:0] SignImmD;

	/*** The following outputs are generated by the Execute pipeline stage ***/

	// The control signal denoting whether a register is written to.
	output reg RegWriteE;

	// The control signal denoting whether data is being written from
	// memory to a register.
	output reg MemtoRegE;

	// The control signal denoting whether main memory is being written to.
	output reg MemWriteE;

	// The four-bit ALU op denoting which operation the ALU should perform.
	output reg [3:0] ALUControlE;

	// The control signal denoting whether the ALU input is an immediate value.
	output reg ALUSrcE;

	// The control signal denoting whether the write reg is rd (R-type instr).
	output reg RegDstE;

	// The data read from the first source register (rs).
	output reg [31:0] RD1E;

	// The data read from the second source register (rt).
	output reg [31:0] RD2E;

	// The first source register.
	output reg [4:0] RsE;

	// The second source register.
	output reg [4:0] RtE;

	// The destination register.
	output reg [4:0] RdE;

	// The sign-extended immediate value.
	output reg [31:0] SignImmE;

	// 1-bit values to propagate
	pipeline_reg_1bit reg_write(clk, FlushE, RegWriteE, RegWriteD);
	pipeline_reg_1bit mem_to_reg(clk, FlushE, MemtoRegE, MemtoRegD);
	pipeline_reg_1bit mem_write(clk, FlushE, MemWriteE, MemWriteD);
	pipeline_reg_1bit alu_src(clk, FlushE, ALUSrcE, ALUSrcD);
	pipeline_reg_1bit reg_dst(clk, FlushE, RegDstE, RegDstD);

	//4-bit values to propagate
	pipeline_reg_4bit alu_control(clk, FlushE, ALUControlE, ALUControlD);

	// 5-bit values to propagate
	pipeline_reg_5bit rs(clk, FlushE, RsE, RsD);
	pipeline_reg_5bit rt(clk, FlushE, RtE, RtD);
	pipeline_reg_5bit rd(clk, FlushE, RdE, RdD);

	// 32-bit values to propagate
	pipeline_reg rd1(clk, FlushE, RD1E, RD1D);
	pipeline_reg rd2(clk, FlushE, RD2E, RD2D);
	pipeline_reg sign_imm(clk, FlushE, SignImmE, SignImmD);

endmodule
`endif

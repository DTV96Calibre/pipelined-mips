`ifndef MIPS_H
`include "mips.h"
`endif

`ifndef MEM_STAGE
`define MEM_STAGE

// This module encapsulates the entire memory pipeline register.
module mem_stage(clk, RegWriteE, MemtoRegE, MemWriteE, ALUOutE, WriteDataE,
	WriteRegE, RegWriteM, MemtoRegM, MemWriteM, ALUOutM, WriteDataM, WriteRegM);

	// The clock.
	input wire clk;

	/*** The following inputs are fed from the Execute pipeline stage ***/

	// The control signal denoting whether a register is written to.
	input wire RegWriteE;

	// The control signal denoting whether data is being written from
	// memory to a register.
	input wire MemtoRegE;

	// The control signal denoting whether main memory is being written to.
	input wire MemWriteE;

	// The 32-bit output computed by the ALU.
	input wire [31:0] ALUOutE;

	// The 32-bit value to write to memory.
	input wire [31:0] WriteDataE;

	// The 5-bit register code that will be written to.
	input wire [4:0] WriteRegE;

	/*** The following outputs are generated by the Memory pipeline stage ***/

	// The control signal denoting whether a register is written to.
	output reg RegWriteM;

	// The control signal denoting whether data is being written from
	// memory to a register.
	output reg MemtoRegM;

	// The control signal denoting whether main memory is being written to.
	output reg MemWriteM;

	// The 32-bit output computed by the ALU.
	output reg [31:0] ALUOutM;

	// The 32-bit value to write to memory.
	output reg [31:0] WriteDataM;

	// The 5-bit register code that will be written to.
	output reg [4:0] WriteRegM;

	// Values in the mem stage will always pass through
	wire signal;
	assign signal = 1;

	// Propagate values
	pipeline_reg_1bit reg_write(clk, signal, RegWriteM, RegWriteE);
	pipeline_reg_1bit mem_to_reg(clk, signal, MemtoRegM, MemtoRegE);
	pipeline_reg_1bit mem_write(clk, signal, MemWriteM, MemWriteE);
	pipeline_reg alu_out(clk, signal, ALUOutM, ALUOutE);
	pipeline_reg write_data(clk, signal, WriteDataM, WriteDataE);
	pipeline_reg_5bit write_reg(clk, signal, WriteRegM, WriteRegE);

endmodule
`endif




`ifndef DECODE_PIPELINE_REG
`define DECODE_PIPELINE_REG

`include "pipeline_reg.v"

module decode_pipeline_reg(clock, 


`endif



